module mem();


reg [7:0] Memory [16'h1000:0];
integer itr;

/*
always @(*)
            begin
            for(ind=0;ind<4;ind=ind+1)
            begin
            Dm1[8*ind +: 8] =  Mem[a1];
            a1 = a1 + 1 ;
            end
            end
*/


endmodule

