`include "vscale_md_constants.vh"
`include "vscale_ctrl_constants.vh"	//Change file name
`include "rv32_opcodes.vh"

`timescale 1ns/1ps

module alu_div_mul(
	input			clk,
	
);